library IEEE;
use IEEE.std_logic_1164.all;

package bullet_tank_const is
    constant bullet_width : integer := 20;
    constant bullet_height : integer := 20;
    constant bullet_speed : integer := 5;

    constant tank_width : integer := 100;
    constant tank_height : integer := 50;

    constant screen_width : integer := 640;
    constant screen_height : integer := 480;
end package bullet_tank_const;
package body bullet_tank_const is
end package body bullet_tank_const;

